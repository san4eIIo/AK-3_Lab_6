library verilog;
use verilog.vl_types.all;
entity lab6v2_vlg_sample_tst is
    port(
        in_x1           : in     vl_logic;
        in_x2           : in     vl_logic;
        in_x3           : in     vl_logic;
        in_x4           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab6v2_vlg_sample_tst;

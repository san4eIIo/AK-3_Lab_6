library verilog;
use verilog.vl_types.all;
entity lab6v2_vlg_check_tst is
    port(
        out_y           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab6v2_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity lab6v2_vlg_vec_tst is
end lab6v2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity lab6v2 is
    port(
        out_y           : out    vl_logic;
        in_x1           : in     vl_logic;
        in_x2           : in     vl_logic;
        in_x3           : in     vl_logic;
        in_x4           : in     vl_logic
    );
end lab6v2;

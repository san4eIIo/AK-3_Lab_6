library verilog;
use verilog.vl_types.all;
entity Lab6_vlg_check_tst is
    port(
        out_y           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab6_vlg_check_tst;
